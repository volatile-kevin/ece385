module registerUnit(
                    input logic [2:0] DR_mux_in,
                    input logic LD.REG,
                    input logic [2:0] SR2,
                    input logic [2:0] SR1_mux_in,
                    input logic [15:0] bus_data,
                    output logic [15:0] SR1_out, SR2_out
);



endmodule