module alu(

);

endmodule